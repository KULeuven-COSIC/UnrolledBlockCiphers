library ieee;
use ieee.std_logic_1164.all;

package constants is
    type round_array is array(5 downto 0) of std_logic_vector(63 downto 0);
end package;
