library ieee;
use ieee.std_logic_1164.all;

entity aes_sbox is
    port (
        datai : in  std_logic_vector(7 downto 0);
        datao : out std_logic_vector(7 downto 0)
    );
end entity;

architecture rtl of aes_sbox is
begin
    lookup_process : process (datai) is
    begin
        lookup_case : case datai is
            when x"00"  => datao <= x"63";
            when x"01"  => datao <= x"7C";
            when x"02"  => datao <= x"77";
            when x"03"  => datao <= x"7B";
            when x"04"  => datao <= x"F2";
            when x"05"  => datao <= x"6B";
            when x"06"  => datao <= x"6F";
            when x"07"  => datao <= x"C5";
            when x"08"  => datao <= x"30";
            when x"09"  => datao <= x"01";
            when x"0A"  => datao <= x"67";
            when x"0B"  => datao <= x"2B";
            when x"0C"  => datao <= x"FE";
            when x"0D"  => datao <= x"D7";
            when x"0E"  => datao <= x"AB";
            when x"0F"  => datao <= x"76";

            when x"10"  => datao <= x"CA";
            when x"11"  => datao <= x"82";
            when x"12"  => datao <= x"C9";
            when x"13"  => datao <= x"7D";
            when x"14"  => datao <= x"FA";
            when x"15"  => datao <= x"59";
            when x"16"  => datao <= x"47";
            when x"17"  => datao <= x"F0";
            when x"18"  => datao <= x"AD";
            when x"19"  => datao <= x"D4";
            when x"1A"  => datao <= x"A2";
            when x"1B"  => datao <= x"AF";
            when x"1C"  => datao <= x"9C";
            when x"1D"  => datao <= x"A4";
            when x"1E"  => datao <= x"72";
            when x"1F"  => datao <= x"C0";

            when x"20"  => datao <= x"B7";
            when x"21"  => datao <= x"FD";
            when x"22"  => datao <= x"93";
            when x"23"  => datao <= x"26";
            when x"24"  => datao <= x"36";
            when x"25"  => datao <= x"3F";
            when x"26"  => datao <= x"F7";
            when x"27"  => datao <= x"CC";
            when x"28"  => datao <= x"34";
            when x"29"  => datao <= x"A5";
            when x"2A"  => datao <= x"E5";
            when x"2B"  => datao <= x"F1";
            when x"2C"  => datao <= x"71";
            when x"2D"  => datao <= x"D8";
            when x"2E"  => datao <= x"31";
            when x"2F"  => datao <= x"15";

            when x"30"  => datao <= x"04";
            when x"31"  => datao <= x"C7";
            when x"32"  => datao <= x"23";
            when x"33"  => datao <= x"C3";
            when x"34"  => datao <= x"18";
            when x"35"  => datao <= x"96";
            when x"36"  => datao <= x"05";
            when x"37"  => datao <= x"9A";
            when x"38"  => datao <= x"07";
            when x"39"  => datao <= x"12";
            when x"3A"  => datao <= x"80";
            when x"3B"  => datao <= x"E2";
            when x"3C"  => datao <= x"EB";
            when x"3D"  => datao <= x"27";
            when x"3E"  => datao <= x"B2";
            when x"3F"  => datao <= x"75";

            when x"40"  => datao <= x"09";
            when x"41"  => datao <= x"83";
            when x"42"  => datao <= x"2C";
            when x"43"  => datao <= x"1A";
            when x"44"  => datao <= x"1B";
            when x"45"  => datao <= x"6E";
            when x"46"  => datao <= x"5A";
            when x"47"  => datao <= x"A0";
            when x"48"  => datao <= x"52";
            when x"49"  => datao <= x"3B";
            when x"4A"  => datao <= x"D6";
            when x"4B"  => datao <= x"B3";
            when x"4C"  => datao <= x"29";
            when x"4D"  => datao <= x"E3";
            when x"4E"  => datao <= x"2F";
            when x"4F"  => datao <= x"84";

            when x"50"  => datao <= x"53";
            when x"51"  => datao <= x"D1";
            when x"52"  => datao <= x"00";
            when x"53"  => datao <= x"ED";
            when x"54"  => datao <= x"20";
            when x"55"  => datao <= x"FC";
            when x"56"  => datao <= x"B1";
            when x"57"  => datao <= x"5B";
            when x"58"  => datao <= x"6A";
            when x"59"  => datao <= x"CB";
            when x"5A"  => datao <= x"BE";
            when x"5B"  => datao <= x"39";
            when x"5C"  => datao <= x"4A";
            when x"5D"  => datao <= x"4C";
            when x"5E"  => datao <= x"58";
            when x"5F"  => datao <= x"CF";

            when x"60"  => datao <= x"D0";
            when x"61"  => datao <= x"EF";
            when x"62"  => datao <= x"AA";
            when x"63"  => datao <= x"FB";
            when x"64"  => datao <= x"43";
            when x"65"  => datao <= x"4D";
            when x"66"  => datao <= x"33";
            when x"67"  => datao <= x"85";
            when x"68"  => datao <= x"45";
            when x"69"  => datao <= x"F9";
            when x"6A"  => datao <= x"02";
            when x"6B"  => datao <= x"7F";
            when x"6C"  => datao <= x"50";
            when x"6D"  => datao <= x"3C";
            when x"6E"  => datao <= x"9F";
            when x"6F"  => datao <= x"A8";

            when x"70"  => datao <= x"51";
            when x"71"  => datao <= x"A3";
            when x"72"  => datao <= x"40";
            when x"73"  => datao <= x"8F";
            when x"74"  => datao <= x"92";
            when x"75"  => datao <= x"9D";
            when x"76"  => datao <= x"38";
            when x"77"  => datao <= x"F5";
            when x"78"  => datao <= x"BC";
            when x"79"  => datao <= x"B6";
            when x"7A"  => datao <= x"DA";
            when x"7B"  => datao <= x"21";
            when x"7C"  => datao <= x"10";
            when x"7D"  => datao <= x"FF";
            when x"7E"  => datao <= x"F3";
            when x"7F"  => datao <= x"D2";

            when x"80"  => datao <= x"CD";
            when x"81"  => datao <= x"0C";
            when x"82"  => datao <= x"13";
            when x"83"  => datao <= x"EC";
            when x"84"  => datao <= x"5F";
            when x"85"  => datao <= x"97";
            when x"86"  => datao <= x"44";
            when x"87"  => datao <= x"17";
            when x"88"  => datao <= x"C4";
            when x"89"  => datao <= x"A7";
            when x"8A"  => datao <= x"7E";
            when x"8B"  => datao <= x"3D";
            when x"8C"  => datao <= x"64";
            when x"8D"  => datao <= x"5D";
            when x"8E"  => datao <= x"19";
            when x"8F"  => datao <= x"73";

            when x"90"  => datao <= x"60";
            when x"91"  => datao <= x"81";
            when x"92"  => datao <= x"4F";
            when x"93"  => datao <= x"DC";
            when x"94"  => datao <= x"22";
            when x"95"  => datao <= x"2A";
            when x"96"  => datao <= x"90";
            when x"97"  => datao <= x"88";
            when x"98"  => datao <= x"46";
            when x"99"  => datao <= x"EE";
            when x"9A"  => datao <= x"B8";
            when x"9B"  => datao <= x"14";
            when x"9C"  => datao <= x"DE";
            when x"9D"  => datao <= x"5E";
            when x"9E"  => datao <= x"0B";
            when x"9F"  => datao <= x"DB";

            when x"A0"  => datao <= x"E0";
            when x"A1"  => datao <= x"32";
            when x"A2"  => datao <= x"3A";
            when x"A3"  => datao <= x"0A";
            when x"A4"  => datao <= x"49";
            when x"A5"  => datao <= x"06";
            when x"A6"  => datao <= x"24";
            when x"A7"  => datao <= x"5C";
            when x"A8"  => datao <= x"C2";
            when x"A9"  => datao <= x"D3";
            when x"AA"  => datao <= x"AC";
            when x"AB"  => datao <= x"62";
            when x"AC"  => datao <= x"91";
            when x"AD"  => datao <= x"95";
            when x"AE"  => datao <= x"E4";
            when x"AF"  => datao <= x"79";

            when x"B0"  => datao <= x"E7";
            when x"B1"  => datao <= x"C8";
            when x"B2"  => datao <= x"37";
            when x"B3"  => datao <= x"6D";
            when x"B4"  => datao <= x"8D";
            when x"B5"  => datao <= x"D5";
            when x"B6"  => datao <= x"4E";
            when x"B7"  => datao <= x"A9";
            when x"B8"  => datao <= x"6C";
            when x"B9"  => datao <= x"56";
            when x"BA"  => datao <= x"F4";
            when x"BB"  => datao <= x"EA";
            when x"BC"  => datao <= x"65";
            when x"BD"  => datao <= x"7A";
            when x"BE"  => datao <= x"AE";
            when x"BF"  => datao <= x"08";

            when x"C0"  => datao <= x"BA";
            when x"C1"  => datao <= x"78";
            when x"C2"  => datao <= x"25";
            when x"C3"  => datao <= x"2E";
            when x"C4"  => datao <= x"1C";
            when x"C5"  => datao <= x"A6";
            when x"C6"  => datao <= x"B4";
            when x"C7"  => datao <= x"C6";
            when x"C8"  => datao <= x"E8";
            when x"C9"  => datao <= x"DD";
            when x"CA"  => datao <= x"74";
            when x"CB"  => datao <= x"1F";
            when x"CC"  => datao <= x"4B";
            when x"CD"  => datao <= x"BD";
            when x"CE"  => datao <= x"8B";
            when x"CF"  => datao <= x"8A";

            when x"D0"  => datao <= x"70";
            when x"D1"  => datao <= x"3E";
            when x"D2"  => datao <= x"B5";
            when x"D3"  => datao <= x"66";
            when x"D4"  => datao <= x"48";
            when x"D5"  => datao <= x"03";
            when x"D6"  => datao <= x"F6";
            when x"D7"  => datao <= x"0E";
            when x"D8"  => datao <= x"61";
            when x"D9"  => datao <= x"35";
            when x"DA"  => datao <= x"57";
            when x"DB"  => datao <= x"B9";
            when x"DC"  => datao <= x"86";
            when x"DD"  => datao <= x"C1";
            when x"DE"  => datao <= x"1D";
            when x"DF"  => datao <= x"9E";

            when x"E0"  => datao <= x"E1";
            when x"E1"  => datao <= x"F8";
            when x"E2"  => datao <= x"98";
            when x"E3"  => datao <= x"11";
            when x"E4"  => datao <= x"69";
            when x"E5"  => datao <= x"D9";
            when x"E6"  => datao <= x"8E";
            when x"E7"  => datao <= x"94";
            when x"E8"  => datao <= x"9B";
            when x"E9"  => datao <= x"1E";
            when x"EA"  => datao <= x"87";
            when x"EB"  => datao <= x"E9";
            when x"EC"  => datao <= x"CE";
            when x"ED"  => datao <= x"55";
            when x"EE"  => datao <= x"28";
            when x"EF"  => datao <= x"DF";
            
            when x"F0"  => datao <= x"8C";
            when x"F1"  => datao <= x"A1";
            when x"F2"  => datao <= x"89";
            when x"F3"  => datao <= x"0D";
            when x"F4"  => datao <= x"BF";
            when x"F5"  => datao <= x"E6";
            when x"F6"  => datao <= x"42";
            when x"F7"  => datao <= x"68";
            when x"F8"  => datao <= x"41";
            when x"F9"  => datao <= x"99";
            when x"FA"  => datao <= x"2D";
            when x"FB"  => datao <= x"0F";
            when x"FC"  => datao <= x"B0";
            when x"FD"  => datao <= x"54";
            when x"FE"  => datao <= x"BB";
            when x"FF"  => datao <= x"16";

            when others => datao <= (others => 'X');
        end case lookup_case;
    end process lookup_process;
end architecture rtl;
